-- Implements a simple Nios II system for the DE2-115 board.
-- Inputs: SW7-0 are parallel port inputs to the Nios II system
-- CLOCK_50 is the system clock
-- KEY0 is the active-low system reset
-- Outputs: LEDG7−0 are parallel port outputs from the Nios II system
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY top_level IS
PORT (
    KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    CLOCK_50 : IN STD_LOGIC;
    LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    UART_TXD : OUT STD_LOGIC;
    UART_RXD : IN STD_LOGIC;
    HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
    HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
    HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
    );
END top_level;

ARCHITECTURE Structure OF top_level IS

component system is
    port (
        clk_clk                         : in  std_logic                    := 'X'; -- clk
        leds_external_connection_export : out std_logic_vector(7 downto 0);        -- export
        reset_reset_n                   : in  std_logic                    := 'X'; -- reset_n
        rs232_0_external_interface_RXD  : in  std_logic                    := 'X'; -- RXD
        rs232_0_external_interface_TXD  : out std_logic;                           -- TXD
        full_display_0_disp0_to_disp    : out std_logic_vector(6 downto 0);        -- to_disp
        full_display_0_disp1_to_disp    : out std_logic_vector(6 downto 0);        -- to_disp
        full_display_0_disp2_to_disp    : out std_logic_vector(6 downto 0)         -- to_disp
    );
end component system;

BEGIN

-- Instantiate the Nios II system entity generated by the SOPC Builder
-- Nios II: nios_system PORT MAP (CLOCK_50, KEY(0), LEDG, SW);
u0 : component system
    port map (
        clk_clk                         => CLOCK_50,                         --                        clk.clk
        leds_external_connection_export => LEDG, --   leds_external_connection.export
        reset_reset_n                   => KEY(0),                   --                      reset.reset_n
        rs232_0_external_interface_RXD  => UART_RXD,  -- rs232_0_external_interface.RXD
        rs232_0_external_interface_TXD  => UART_TXD,  --                           .TXD
        full_display_0_disp0_to_disp    => HEX0,    --       full_display_0_disp0.to_disp
        full_display_0_disp1_to_disp    => HEX1,    --       full_display_0_disp1.to_disp
        full_display_0_disp2_to_disp    => HEX2     --       full_display_0_disp2.to_disp
    );

END Structure;