-- Implements a simple Nios II system for the DE2-115 board.
-- Inputs: SW7-0 are parallel port inputs to the Nios II system
-- CLOCK_50 is the system clock
-- KEY0 is the active-low system reset
-- Outputs: LEDG7−0 are parallel port outputs from the Nios II system
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY top_level IS
PORT (
    -- Add all required ports here, their names should match what is in 'DE2_115_pin_assignments.csv'
    KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    CLOCK_50 : IN STD_LOGIC;
    LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    UART_TXD : OUT STD_LOGIC;
    UART_RXD : IN STD_LOGIC
    );
END top_level;

ARCHITECTURE Structure OF top_level IS

-- Copy the system component declaration here from system_inst.vhd
component system is
    port (
        clk_clk                         : in  std_logic                    := 'X'; -- clk
        reset_reset_n                   : in  std_logic                    := 'X'; -- reset_n
        rs232_0_external_interface_RXD  : in  std_logic                    := 'X'; -- RXD
        rs232_0_external_interface_TXD  : out std_logic;                           -- TXD
        leds_external_connection_export : out std_logic_vector(7 downto 0)         -- export
    );
end component system;

BEGIN

-- Instantiate the Nios II system entity generated by the SOPC Builder and connect it to the pins
u0 : component system
    port map (
        clk_clk                         => CLOCK_50,        --                        clk.clk
        reset_reset_n                   => KEY(0),          --                      reset.reset_n
        rs232_0_external_interface_RXD  => UART_RXD,        -- rs232_0_external_interface.RXD
        rs232_0_external_interface_TXD  => UART_TXD,        --                           .TXD
        leds_external_connection_export => LEDG             --   leds_external_connection.export
    );

END Structure;